library ieee;
use ieee.std_logic_1164.all;


entity InfraredReciver is
	port (
		clk : in std_logic;
		rst : in std_logic
	);
end entity InfraredReciver;

architecture InfraredReciver_Arc of InfraredReciver is
	
begin

	
end architecture InfraredReciver_Arc;