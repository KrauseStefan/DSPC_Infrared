library ieee;
use ieee.std_logic_1164.all;

-------------------------------------------------------------------------------

entity IF_Receiver_TB is
  
end IF_Receiver_TB;

-------------------------------------------------------------------------------

architecture test of IF_Receiver_TB is

begin
  
end test;