
library ieee;
use ieee.std_logic_1164.all;

entity Counter is
	port (
		clk : in std_logic;
		rst : in std_logic
	);
end entity Counter;
