library ieee;
use ieee.std_logic_1164.all;


entity BitSampler is
	port (
		clk : in std_logic;
		rst : in std_logic
	);
end entity BitSampler;


architecture BitSamplerArc of BitSampler is
	
begin
	
end architecture BitSamplerArc;